`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:43:01 12/25/2013 
// Design Name: 
// Module Name:    alu 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module alu (alu_zero_flag, alu_out, data_1, data_2, sel);
  
	// Opcodes
	wire [`WORD_SIZE:0] sub_res;
	wire [`WORD_SIZE:0] add_res;
	
	wire oflow_add;	//�ӷ����λ
	wire oflow_sub;	//�������λ 
	wire oflow;			//�ܵ����λ
	
	output alu_zero_flag;
	output [`WORD_SIZE-1: 0] alu_out;
	input [`WORD_SIZE-1: 0] data_1, data_2;
	input [`OP_SIZE-1: 0] sel;
	
	assign sub_res = data_1 - data_2;
	assign add_res = data_1 + data_2;
	
	assign oflow_sub = (data_1[`WORD_SIZE-1] != data_2[`WORD_SIZE-1] && sub_res[`WORD_SIZE-1] == data_2[`WORD_SIZE-1]) ? 1 : 0;
	assign oflow_add = (data_1[`WORD_SIZE-1] == data_2[`WORD_SIZE-1] && add_res[`WORD_SIZE-1] != data_1[`WORD_SIZE-1]) ? 1 : 0;
  
	reg [`WORD_SIZE-1: 0] 	alu_out;
	assign  alu_zero_flag = (0 == alu_out);
	always @ (*)  
		case  (sel)
			`ADD: alu_out <= add_res;
			`OR: alu_out <= data_1 | data_2;
			`SUB: alu_out <= sub_res;
			`AND: alu_out <= data_1 & data_2;
			`SLT: alu_out <= (data_1 < data_2) ? 1: 0;
			default: alu_out <= 0;
		endcase 
endmodule
